
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY SumadorTB IS
END SumadorTB;
 
ARCHITECTURE behavior OF SumadorTB IS 
 
 
    COMPONENT Sumador
    PORT(
         In1 : IN  std_logic_vector(31 downto 0);
         In2 : IN  std_logic_vector(31 downto 0);
         Out1 : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal In1 : std_logic_vector(31 downto 0) := (others => '0');
   signal In2 : std_logic_vector(31 downto 0) := (others => '0');

 	--Outputs
   signal Out1 : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Sumador PORT MAP (
          In1 => In1,
          In2 => In2,
          Out1 => Out1
        );
 

   -- Stimulus process
   stim_proc: process
   begin
	Out1<= In1+In2;
	

      wait;
   end process;

END;
