----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:24:24 10/06/2017 
-- Design Name: 
-- Module Name:    Mux1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Mux1 is
    Port ( In1 : in  STD_LOGIC_VECTOR (31 downto 0);
           In2 : in  STD_LOGIC_VECTOR (31 downto 0);
           i : in  STD_LOGIC;
           outMux : out STD_LOGIC_VECTOR (31 downto 0));
end Mux1;

architecture Behavioral of Mux1 is

begin
process(In1,In2,i)
       begin 
		  
		  case i is 
		     
			  when '0' => 
			  outMux <= In1;
			  
			  when '1' =>
			  outMux <= In2;
			  
			  when others =>
			  outMux <= "00000000000000000000000000000000";

        end case;
end process;
end Behavioral;

